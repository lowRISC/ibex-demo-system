../../../../ibex-demo-system-labs/lab4_supplementary_material/fp_mul.sv